library verilog;
use verilog.vl_types.all;
entity cc_1 is
    port(
        rst             : in     vl_logic;
        start           : in     vl_logic;
        m0              : in     vl_logic_vector(15 downto 0);
        m1              : in     vl_logic_vector(15 downto 0);
        clk             : in     vl_logic;
        index           : out    vl_logic_vector(15 downto 0);
        done            : out    vl_logic
    );
end cc_1;
